// MUX

module VGAmux (


); 



endmodule