/*
Vending Machine Top with FSM 
*/ 