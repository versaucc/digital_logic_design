// Decoder

module VGAdecoder (

);


endmodule